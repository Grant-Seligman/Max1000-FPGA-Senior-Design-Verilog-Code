// adc_core.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module adc_core (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         pll_c0_clk;                                       // pll:c0 -> adc:adc_pll_clock_clk
	wire         pll_locked_conduit_export;                        // pll:locked -> adc:adc_pll_locked_export
	wire  [31:0] avalon_bridge_master_readdata;                    // mm_interconnect_0:avalon_bridge_master_readdata -> avalon_bridge:master_readdata
	wire         avalon_bridge_master_waitrequest;                 // mm_interconnect_0:avalon_bridge_master_waitrequest -> avalon_bridge:master_waitrequest
	wire  [31:0] avalon_bridge_master_address;                     // avalon_bridge:master_address -> mm_interconnect_0:avalon_bridge_master_address
	wire         avalon_bridge_master_read;                        // avalon_bridge:master_read -> mm_interconnect_0:avalon_bridge_master_read
	wire   [3:0] avalon_bridge_master_byteenable;                  // avalon_bridge:master_byteenable -> mm_interconnect_0:avalon_bridge_master_byteenable
	wire         avalon_bridge_master_readdatavalid;               // mm_interconnect_0:avalon_bridge_master_readdatavalid -> avalon_bridge:master_readdatavalid
	wire         avalon_bridge_master_write;                       // avalon_bridge:master_write -> mm_interconnect_0:avalon_bridge_master_write
	wire  [31:0] avalon_bridge_master_writedata;                   // avalon_bridge:master_writedata -> mm_interconnect_0:avalon_bridge_master_writedata
	wire  [31:0] mm_interconnect_0_adc_sample_store_csr_readdata;  // adc:sample_store_csr_readdata -> mm_interconnect_0:adc_sample_store_csr_readdata
	wire   [6:0] mm_interconnect_0_adc_sample_store_csr_address;   // mm_interconnect_0:adc_sample_store_csr_address -> adc:sample_store_csr_address
	wire         mm_interconnect_0_adc_sample_store_csr_read;      // mm_interconnect_0:adc_sample_store_csr_read -> adc:sample_store_csr_read
	wire         mm_interconnect_0_adc_sample_store_csr_write;     // mm_interconnect_0:adc_sample_store_csr_write -> adc:sample_store_csr_write
	wire  [31:0] mm_interconnect_0_adc_sample_store_csr_writedata; // mm_interconnect_0:adc_sample_store_csr_writedata -> adc:sample_store_csr_writedata
	wire  [31:0] mm_interconnect_0_adc_sequencer_csr_readdata;     // adc:sequencer_csr_readdata -> mm_interconnect_0:adc_sequencer_csr_readdata
	wire   [0:0] mm_interconnect_0_adc_sequencer_csr_address;      // mm_interconnect_0:adc_sequencer_csr_address -> adc:sequencer_csr_address
	wire         mm_interconnect_0_adc_sequencer_csr_read;         // mm_interconnect_0:adc_sequencer_csr_read -> adc:sequencer_csr_read
	wire         mm_interconnect_0_adc_sequencer_csr_write;        // mm_interconnect_0:adc_sequencer_csr_write -> adc:sequencer_csr_write
	wire  [31:0] mm_interconnect_0_adc_sequencer_csr_writedata;    // mm_interconnect_0:adc_sequencer_csr_writedata -> adc:sequencer_csr_writedata
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [adc:reset_sink_reset_n, mm_interconnect_0:adc_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_0:avalon_bridge_clk_reset_reset_bridge_in_reset_reset, pll:reset]

	adc_core_adc adc (
		.clock_clk                  (clk_clk),                                          //            clock.clk
		.reset_sink_reset_n         (~rst_controller_reset_out_reset),                  //       reset_sink.reset_n
		.adc_pll_clock_clk          (pll_c0_clk),                                       //    adc_pll_clock.clk
		.adc_pll_locked_export      (pll_locked_conduit_export),                        //   adc_pll_locked.export
		.sequencer_csr_address      (mm_interconnect_0_adc_sequencer_csr_address),      //    sequencer_csr.address
		.sequencer_csr_read         (mm_interconnect_0_adc_sequencer_csr_read),         //                 .read
		.sequencer_csr_write        (mm_interconnect_0_adc_sequencer_csr_write),        //                 .write
		.sequencer_csr_writedata    (mm_interconnect_0_adc_sequencer_csr_writedata),    //                 .writedata
		.sequencer_csr_readdata     (mm_interconnect_0_adc_sequencer_csr_readdata),     //                 .readdata
		.sample_store_csr_address   (mm_interconnect_0_adc_sample_store_csr_address),   // sample_store_csr.address
		.sample_store_csr_read      (mm_interconnect_0_adc_sample_store_csr_read),      //                 .read
		.sample_store_csr_write     (mm_interconnect_0_adc_sample_store_csr_write),     //                 .write
		.sample_store_csr_writedata (mm_interconnect_0_adc_sample_store_csr_writedata), //                 .writedata
		.sample_store_csr_readdata  (mm_interconnect_0_adc_sample_store_csr_readdata),  //                 .readdata
		.sample_store_irq_irq       ()                                                  // sample_store_irq.irq
	);

	adc_core_avalon_bridge #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) avalon_bridge (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                     //    clk_reset.reset
		.master_address       (avalon_bridge_master_address),       //       master.address
		.master_readdata      (avalon_bridge_master_readdata),      //             .readdata
		.master_read          (avalon_bridge_master_read),          //             .read
		.master_write         (avalon_bridge_master_write),         //             .write
		.master_writedata     (avalon_bridge_master_writedata),     //             .writedata
		.master_waitrequest   (avalon_bridge_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (avalon_bridge_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (avalon_bridge_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	adc_core_pll pll (
		.clk                (clk_clk),                        //       inclk_interface.clk
		.reset              (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read               (),                               //             pll_slave.read
		.write              (),                               //                      .write
		.address            (),                               //                      .address
		.readdata           (),                               //                      .readdata
		.writedata          (),                               //                      .writedata
		.c0                 (pll_c0_clk),                     //                    c0.clk
		.areset             (),                               //        areset_conduit.export
		.locked             (pll_locked_conduit_export),      //        locked_conduit.export
		.scandone           (),                               //           (terminated)
		.scandataout        (),                               //           (terminated)
		.c1                 (),                               //           (terminated)
		.c2                 (),                               //           (terminated)
		.c3                 (),                               //           (terminated)
		.c4                 (),                               //           (terminated)
		.phasedone          (),                               //           (terminated)
		.phasecounterselect (3'b000),                         //           (terminated)
		.phaseupdown        (1'b0),                           //           (terminated)
		.phasestep          (1'b0),                           //           (terminated)
		.scanclk            (1'b0),                           //           (terminated)
		.scanclkena         (1'b0),                           //           (terminated)
		.scandata           (1'b0),                           //           (terminated)
		.configupdate       (1'b0)                            //           (terminated)
	);

	adc_core_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                       (clk_clk),                                          //                                     clk_0_clk.clk
		.adc_reset_sink_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                   //          adc_reset_sink_reset_bridge_in_reset.reset
		.avalon_bridge_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // avalon_bridge_clk_reset_reset_bridge_in_reset.reset
		.avalon_bridge_master_address                        (avalon_bridge_master_address),                     //                          avalon_bridge_master.address
		.avalon_bridge_master_waitrequest                    (avalon_bridge_master_waitrequest),                 //                                              .waitrequest
		.avalon_bridge_master_byteenable                     (avalon_bridge_master_byteenable),                  //                                              .byteenable
		.avalon_bridge_master_read                           (avalon_bridge_master_read),                        //                                              .read
		.avalon_bridge_master_readdata                       (avalon_bridge_master_readdata),                    //                                              .readdata
		.avalon_bridge_master_readdatavalid                  (avalon_bridge_master_readdatavalid),               //                                              .readdatavalid
		.avalon_bridge_master_write                          (avalon_bridge_master_write),                       //                                              .write
		.avalon_bridge_master_writedata                      (avalon_bridge_master_writedata),                   //                                              .writedata
		.adc_sample_store_csr_address                        (mm_interconnect_0_adc_sample_store_csr_address),   //                          adc_sample_store_csr.address
		.adc_sample_store_csr_write                          (mm_interconnect_0_adc_sample_store_csr_write),     //                                              .write
		.adc_sample_store_csr_read                           (mm_interconnect_0_adc_sample_store_csr_read),      //                                              .read
		.adc_sample_store_csr_readdata                       (mm_interconnect_0_adc_sample_store_csr_readdata),  //                                              .readdata
		.adc_sample_store_csr_writedata                      (mm_interconnect_0_adc_sample_store_csr_writedata), //                                              .writedata
		.adc_sequencer_csr_address                           (mm_interconnect_0_adc_sequencer_csr_address),      //                             adc_sequencer_csr.address
		.adc_sequencer_csr_write                             (mm_interconnect_0_adc_sequencer_csr_write),        //                                              .write
		.adc_sequencer_csr_read                              (mm_interconnect_0_adc_sequencer_csr_read),         //                                              .read
		.adc_sequencer_csr_readdata                          (mm_interconnect_0_adc_sequencer_csr_readdata),     //                                              .readdata
		.adc_sequencer_csr_writedata                         (mm_interconnect_0_adc_sequencer_csr_writedata)     //                                              .writedata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
