
module nios_sys (
	byte_pio_export,
	clk_clk,
	reset_reset_n);	

	output	[3:0]	byte_pio_export;
	input		clk_clk;
	input		reset_reset_n;
endmodule
