
module nios_sys (
	clk_clk,
	reset_reset_n,
	pio_data_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[3:0]	pio_data_export;
endmodule
