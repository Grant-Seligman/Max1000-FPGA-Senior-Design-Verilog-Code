
module nios_sys (
	clk_clk,
	pio_byte_display_export,
	reset_reset_n);	

	input		clk_clk;
	output	[7:0]	pio_byte_display_export;
	input		reset_reset_n;
endmodule
