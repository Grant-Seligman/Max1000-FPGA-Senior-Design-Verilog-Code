
module nios_sys (
	clk_clk,
	reset_reset_n,
	pio_pwm_data_export);	

	input		clk_clk;
	input		reset_reset_n;
	output	[7:0]	pio_pwm_data_export;
endmodule
